`include "base_test.sv"

`include "seq_i2c.sv"

`include "test_dummy.sv"

`include "seq_clk.sv"

`include "test_def_values.sv"

`include "random_test_def_values.sv"

`include "test_w_r_permissions.sv"
